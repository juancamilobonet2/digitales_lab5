/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module CC_COMPARATOR (
//////////// OUTPUTS //////////
	CC_COMPARATOR_result_Out,
//////////// INPUTS //////////
	CC_COMPARATOR_c0_InBUS, // ADDER out
	CC_COMPARATOR_c1_InBUS  // theta
);
//=======================================================
//  PARAMETER declarations
//=======================================================
parameter NUMBER_DATAWIDTH = 8;
//=======================================================
//  PORT declarations
//=======================================================
output reg CC_COMPARATOR_result_Out;
input 	[NUMBER_DATAWIDTH-1:0] CC_COMPARATOR_c0_InBUS;
input 	[NUMBER_DATAWIDTH-1:0] CC_COMPARATOR_c1_InBUS;
//=======================================================
//  REG/WIRE declarations
//=======================================================

//=======================================================
//  Structural coding
//=======================================================
always @(*)
	if (CC_COMPARATOR_c0_InBUS >= CC_COMPARATOR_c1_InBUS)
		CC_COMPARATOR_result_Out=1;
	else
		CC_COMPARATOR_result_Out=0;

endmodule

